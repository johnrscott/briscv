module instr_fetch_unit(
   axi4_lite_if.manager imem_bus
);

   
endmodule
